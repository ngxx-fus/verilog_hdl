module and(
    input A,
    input B,
    input Y
);
    assign Y = A&B;
endmodule