module not (
    input A,
    output Y,
);
    assign y = ~A;
endmodule