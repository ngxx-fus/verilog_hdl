module BIN2BCD(
    input [6:0] BIN,
    output [7:0] BCD
);
    assign BCD = (BIN==0)?(8'H00):(BIN==1)?(8'H01):
    (BIN==2)?(8'H02):(BIN==3)?(8'H03):(BIN==4)?(8'H04):
    (BIN==5)?(8'H05):(BIN==6)?(8'H06):(BIN==7)?(8'H07):
    (BIN==8)?(8'H08):(BIN==9)?(8'H09):(BIN==10)?(8'H10):
    (BIN==11)?(8'H11):(BIN==12)?(8'H12):(BIN==13)?(8'H13):
    (BIN==14)?(8'H14):(BIN==15)?(8'H15):(BIN==16)?(8'H16):
    (BIN==17)?(8'H17):(BIN==18)?(8'H18):(BIN==19)?(8'H19):
    (BIN==20)?(8'H20):(BIN==21)?(8'H21):(BIN==22)?(8'H22):
    (BIN==23)?(8'H23):(BIN==24)?(8'H24):(BIN==25)?(8'H25):
    (BIN==26)?(8'H26):(BIN==27)?(8'H27):(BIN==28)?(8'H28):
    (BIN==29)?(8'H29):
    (BIN==30)?(8'H30):(BIN==31)?(8'H31):(BIN==32)?(8'H32):
    (BIN==33)?(8'H33):(BIN==34)?(8'H34):(BIN==35)?(8'H35):
    (BIN==36)?(8'H36):(BIN==37)?(8'H37):(BIN==38)?(8'H38):
    (BIN==39)?(8'H39):(BIN==40)?(8'H40):(BIN==41)?(8'H41):
    (BIN==42)?(8'H42):(BIN==43)?(8'H43):(BIN==44)?(8'H44):
    (BIN==45)?(8'H45):(BIN==46)?(8'H46):(BIN==47)?(8'H47):
    (BIN==48)?(8'H48):(BIN==49)?(8'H49):(BIN==50)?(8'H50):
    (BIN==51)?(8'H51):(BIN==52)?(8'H52):(BIN==53)?(8'H53):
    (BIN==54)?(8'H54):(BIN==55)?(8'H55):(BIN==56)?(8'H56):
    (BIN==57)?(8'H57):(BIN==58)?(8'H58):(BIN==59)?(8'H59):
    (BIN==60)?(8'H60):(BIN==61)?(8'H61):(BIN==62)?(8'H62):
    (BIN==63)?(8'H63):(BIN==64)?(8'H64):(BIN==65)?(8'H65):
    (BIN==66)?(8'H66):(BIN==67)?(8'H67):(BIN==68)?(8'H68):
    (BIN==69)?(8'H69):(BIN==70)?(8'H70):(BIN==71)?(8'H71):
    (BIN==72)?(8'H72):(BIN==73)?(8'H73):(BIN==74)?(8'H74):
    (BIN==75)?(8'H75):(BIN==76)?(8'H76):(BIN==77)?(8'H77):
    (BIN==78)?(8'H78):(BIN==79)?(8'H79):(BIN==80)?(8'H80):
    (BIN==81)?(8'H81):(BIN==82)?(8'H82):(BIN==83)?(8'H83):
    (BIN==84)?(8'H84):(BIN==85)?(8'H85):(BIN==86)?(8'H86):
    (BIN==87)?(8'H87):(BIN==88)?(8'H88):(BIN==89)?(8'H89):
    (BIN==90)?(8'H90):(BIN==91)?(8'H91):(BIN==92)?(8'H92):
    (BIN==93)?(8'H93):(BIN==94)?(8'H94):(BIN==95)?(8'H95):
    (BIN==96)?(8'H96):(BIN==97)?(8'H97):(BIN==98)?(8'H98):
    (BIN==99)?(8'H99):(8'H99);

endmodule